library IEEE;
library work;
use work.custom_types.all;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Controller_tb is
--  Port ( );
end Controller_tb;

architecture Behavioral of Controller_tb is


component Controller is
    Port (
        ------------------------------------------------  
        ------------------------------------------------  
        -- INPUTS
        clk_in:in STD_LOGIC;
        rst: in STD_LOGIC;
        incoming_inst: in STD_LOGIC;   
        ------------------------------------------------  
        vect_inst : in STD_LOGIC_VECTOR (31 downto 0);
        
        CSR_Addr: in STD_LOGIC_VECTOR ( 11 downto 0);   -- reg address of the CSR                 -- 11 is based on spec sheet
        CSR_WD: in STD_LOGIC_VECTOR (XLEN-1 downto 0); 
        CSR_WEN: in STD_LOGIC;
        rs1_data: in STD_LOGIC_VECTOR( XLEN-1 downto 0);  
        rs2_data: in STD_LOGIC_VECTOR(XLEN-1 downto 0);
        i_done: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --done flag generated by offset_gen and coming from WB pipeline reg (to align with end of write/end of instruction) 
        ------------------------------------------------   
        ------------------------------------------------      
        -- OUTPUTS  
        rd_data: out STD_LOGIC_VECTOR (XLEN-1 downto 0);  --to scalar slave register  
        WriteEn : out STD_LOGIC_VECTOR(NB_LANES-1 downto 0); -- enables write to the reg file
        SrcB : out STD_LOGIC_VECTOR(2*NB_LANES-1 downto 0); -- selects between scalar/vector reg or immediate
                                                    -- 00 = vector reg
                                                    -- 01 = scalar reg
                                                    -- 10 = immediate
                                                    -- 11 = RESERVED
        MemWrite : out STD_LOGIC_VECTOR(NB_LANES-1 downto 0);                -- enables write to memory
        MemRead: out STD_LOGIC_VECTOR(NB_LANES-1 downto 0);                  -- enables read from memory
        WBSrc : out STD_LOGIC_VECTOR(NB_LANES-1 downto 0);                    -- selects if wrbsc is from ALU or mem 
                                                    -- 0 = ALU
                                                    -- 1 = Mem    
        CSR_out: out STD_LOGIC_VECTOR (XLEN-1 downto 0);
        ---- 1) vtype fields:
        vill: out STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
        vma:out STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
        vta:out STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
        vlmul: out STD_LOGIC_VECTOR(3*NB_LANES-1 downto 0);  
        sew: out STD_LOGIC_VECTOR (3*NB_LANES-1 downto 0);
        vstart: out STD_LOGIC_VECTOR(lgVLEN*NB_LANES-1 downto 0);
        vl: out STD_LOGIC_VECTOR(XLEN*NB_LANES-1 downto 0);      
        ------------------------------------------------------------------------
        funct6 : out STD_LOGIC_VECTOR (6*NB_LANES-1 downto 0);
        nf : out STD_LOGIC_VECTOR (3*NB_LANES-1 downto 0);
        mop: out STD_LOGIC_VECTOR (2*NB_LANES-1 downto 0);-- goes to memory lane
                                                              -- 00 if unit stride    
                                                              -- 01 reserved
                                                              -- 10 if strided 
                                                              -- 11 if indexed 
        vm : out STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
        vs2_rs2 : out STD_LOGIC_VECTOR (4*NB_LANES-1 downto 0); -- 2nd vector operand
        rs1 : out STD_LOGIC_VECTOR (4*NB_LANES-1 downto 0); --1st vector operand
        RegSel: out STD_LOGIC_VECTOR((READ_PORTS_PER_LANE*NB_LANES*REGS_PER_BANK)-1 downto 0); --going to RegFile_ALU
        WriteDest : out STD_LOGIC_VECTOR (NB_LANES*REGS_PER_BANK-1 downto 0);--going to RegFile_ALU
        Xdata_in: in STD_LOGIC_VECTOR(XLEN-1 downto 0); --data coming from scalar register
        Xdata: out STD_LOGIC_VECTOR(NB_LANES*XLEN-1 downto 0); --data from scalar register, going to RegFile_ALU
        Idata: out STD_LOGIC_VECTOR(NB_LANES*5-1 downto 0); --data coming from immediate field of size 5 bits, going to RegFile_ALU
        funct3_width : out STD_LOGIC_VECTOR (3*NB_LANES-1 downto 0);
        vd_vs3 : out STD_LOGIC_VECTOR (4*NB_LANES-1 downto 0); --vector write destination  
        extension: out STD_LOGIC_VECTOR(NB_LANES-1 downto 0);        -- goes to memory
                                                                     -- 0 if zero extended
                                                                     -- 1 if sign extended    
        memwidth: out STD_LOGIC_VECTOR(4*NB_LANES-1 downto 0);   -- goes to memory,FOLLOWS CUSTOM ENCODING: represents the exponent of the memory element width 
                                                                 -- number of bits/transfer 
        newInst_out: out STD_LOGIC_VECTOR(NB_LANES-1 downto 0)                                             
    );
end component;


signal  clk_in: STD_LOGIC;
signal  rst:  STD_LOGIC;
signal  incoming_inst:  STD_LOGIC;   
signal  CSR_Addr:  STD_LOGIC_VECTOR ( 11 downto 0);   -- reg address of the CSR                 -- 11 is based on spec sheet
signal  CSR_WD:  STD_LOGIC_VECTOR (XLEN-1 downto 0); 
signal  CSR_WEN:  STD_LOGIC;
signal  rs1_data:  STD_LOGIC_VECTOR( XLEN-1 downto 0);  
signal  rs2_data:  STD_LOGIC_VECTOR(XLEN-1 downto 0);
signal  i_done:  STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --done flag generated by offset_gen and coming from WB pipeline reg (to align with end of write/end of instruction) 
signal  rd_data:  STD_LOGIC_VECTOR (XLEN-1 downto 0);  --to scalar slave register  
signal  WriteEn :  STD_LOGIC_VECTOR(NB_LANES-1 downto 0); -- enables write to the reg file
signal  SrcB :  STD_LOGIC_VECTOR(2*NB_LANES-1 downto 0); -- selects between scalar/vector reg or immediate
signal  MemWrite :  STD_LOGIC_VECTOR(NB_LANES-1 downto 0);                -- enables write to memory
signal  MemRead:  STD_LOGIC_VECTOR(NB_LANES-1 downto 0);                  -- enables read from memory
signal  WBSrc :  STD_LOGIC_VECTOR(NB_LANES-1 downto 0);                    -- selects if wrbsc is from ALU or mem 
signal  CSR_out:  STD_LOGIC_VECTOR (XLEN-1 downto 0);
signal  vill:  STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
signal  vma: STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
signal  vta: STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
signal  vlmul:  STD_LOGIC_VECTOR(3*NB_LANES-1 downto 0);  
signal  sew:  STD_LOGIC_VECTOR (3*NB_LANES-1 downto 0);
signal  vstart:  STD_LOGIC_VECTOR(lgVLEN*NB_LANES-1 downto 0);
signal  vl:  STD_LOGIC_VECTOR(XLEN*NB_LANES-1 downto 0);      
signal  funct6 :  STD_LOGIC_VECTOR (6*NB_LANES-1 downto 0);
signal  nf :  STD_LOGIC_VECTOR (3*NB_LANES-1 downto 0);
signal  mop:  STD_LOGIC_VECTOR (2*NB_LANES-1 downto 0);-- goes to memory lane
signal  vm :  STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
signal  vs2_rs2 :  STD_LOGIC_VECTOR (4*NB_LANES-1 downto 0); -- 2nd vector operand
signal  rs1 :  STD_LOGIC_VECTOR (4*NB_LANES-1 downto 0); --1st vector operand
signal  RegSel:  STD_LOGIC_VECTOR((READ_PORTS_PER_LANE*NB_LANES*REGS_PER_BANK)-1 downto 0); --going to RegFile_ALU
signal  WriteDest :  STD_LOGIC_VECTOR (NB_LANES*REGS_PER_BANK-1 downto 0);--going to RegFile_ALU
signal  Xdata_in:  STD_LOGIC_VECTOR(XLEN-1 downto 0); --data coming from scalar register
signal  Xdata:  STD_LOGIC_VECTOR(NB_LANES*XLEN-1 downto 0); --data from scalar register, going to RegFile_ALU
signal  Idata:  STD_LOGIC_VECTOR(NB_LANES*5-1 downto 0); --data coming from immediate field of size 5 bits, going to RegFile_ALU
signal  funct3_width :  STD_LOGIC_VECTOR (3*NB_LANES-1 downto 0);
signal  vd_vs3 :  STD_LOGIC_VECTOR (4*NB_LANES-1 downto 0); --vector write destination  
signal  extension:  STD_LOGIC_VECTOR(NB_LANES-1 downto 0);        -- goes to memory
signal  memwidth:  STD_LOGIC_VECTOR(4*NB_LANES-1 downto 0);   -- goes to memory,FOLLOWS CUSTOM ENCODING: represents the exponent of the memory element width 
signal  newInst_out:  STD_LOGIC_VECTOR(NB_LANES-1 downto 0);



-- The following signals are used to make testing each instruction easier
signal    t_vect_inst: STD_LOGIC_VECTOR(31 downto 0); 
signal    t_vs1: STD_LOGIC_VECTOR(4 downto 0);
signal    t_vs2: STD_LOGIC_VECTOR(4 downto 0);
signal    t_vd: STD_LOGIC_VECTOR(4 downto 0);
signal    t_opcode: STD_LOGIC_VECTOR(6 downto 0);
signal    t_funct3: STD_LOGIC_VECTOR(2 downto 0);
signal    t_funct6: STD_LOGIC_VECTOR(5 downto 0);
signal    t_vm: STD_LOGIC;

begin
t_vect_inst<= t_funct6 & t_vm & t_vs2 & t_vs1 & t_funct3 & t_vd & t_opcode;
    G1: Controller
--    GENERIC MAP(NB_LANES,lgNB_LANES,READ_PORTS_PER_LANE,REGS_PER_BANK,XLEN,VLEN,ELEN,lgELEN,lgVLEN)
    PORT MAP(
            clk_in        =>clk_in        ,
            rst           =>rst           ,
            incoming_inst =>incoming_inst ,
            vect_inst     =>t_vect_inst     ,
            CSR_Addr      =>CSR_Addr      ,
            CSR_WD        =>CSR_WD        ,
            CSR_WEN       =>CSR_WEN       ,
            rs1_data      =>rs1_data      ,
            rs2_data      =>rs2_data      ,
            i_done        =>i_done        ,
            rd_data       =>rd_data       ,
            WriteEn       =>WriteEn       ,
            SrcB          =>SrcB          ,
            MemWrite      =>MemWrite      ,
            MemRead       =>MemRead       ,
            WBSrc         =>WBSrc         ,
            CSR_out       =>CSR_out       ,
            vill          =>vill          ,
            vma           =>vma           ,
            vta           =>vta           ,
            vlmul         =>vlmul         ,
            sew           =>sew           ,
            vstart        =>vstart        ,
            vl            =>vl            ,
            funct6        =>funct6        ,
            nf            =>nf            ,
            mop           =>mop           ,
            vm            =>vm            ,
            vs2_rs2       =>vs2_rs2       ,
            rs1           =>rs1           ,
            RegSel        =>RegSel        ,
            WriteDest     =>WriteDest     ,
            Xdata_in      =>Xdata_in      ,
            Xdata         =>Xdata         ,
            Idata         =>Idata         ,
            funct3_width  =>funct3_width  ,
            vd_vs3        =>vd_vs3        ,
--            extension     =>extension     ,
--            memwidth      =>memwidth      ,
            newInst_out   =>newInst_out   
     );
     
    clk_proc: process begin
        clk_in<='0';
        wait for 5ns;
        clk_in<='1'; 
        wait for 5ns;
    end process;

    process begin
        incoming_inst<='0';rst<='1'; wait for 5 ns; rst<='0'; wait for 5ns;rst<='1';wait for 5 ns;
        --set vstart as 0
        CSR_Addr<=x"008"; CSR_WD<=x"00000000"; CSR_WEN<='1'; wait for 10ns;
        CSR_WEN<='0';
        --vsetvli configuration instruction
        incoming_inst<='1';
        t_funct6<="000000";t_vm<='0';t_vs2<="00000";t_vs1<="00000";t_funct3<="111";t_vd<="00001";t_opcode<="1010111";
        wait for 10 ns;
        incoming_inst<='0';
        wait for 10ns;
--        -- move instruction to fill v0 register
        incoming_inst<='1'; 
        Xdata_in<=x"00000001";
        t_funct6<="010111";t_vm<='1';t_vs2<="00000";t_vs1<="00000";t_funct3<="100";t_vd<="00000";t_opcode<="1010111";
        wait for 10 ns; incoming_inst<='0';  
        wait for 10ns; 
        --move instruction to fill v16 register
        incoming_inst<='1'; 
        Xdata_in<=x"00000002";
        t_funct6<="010111";t_vm<='1';t_vs2<="10100";t_vs1<="10000";t_funct3<="100";t_vd<="10000";t_opcode<="1010111";
        wait for 10 ns; incoming_inst<='0';
        wait for 10ns; 
        -- add immediate instruction on lane 1; adds 4 to v0, and writes sum in v2
        incoming_inst<='1';
        t_funct6<="000000";t_vm<='1';t_vs2<="00000";t_vs1<="00100";t_funct3<="011";t_vd<="00010";t_opcode<="1010111";
        wait for 10 ns; incoming_inst<='0';   
        
        wait;
    end process;

end Behavioral;
