library IEEE;
library work;
use work.custom_types.all;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ALU_with_pipeline_tb is
end ALU_with_pipeline_tb;

architecture ALU_with_pipeline_tb_arch of ALU_with_pipeline_tb is

component ALU_with_pipeline is
    Port (  clk: in STD_LOGIC; 
            rst: in STD_LOGIC;
            mask_reg: in STD_LOGIC_VECTOR(VLEN-1 downto 0);
            vm: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
            sew: in STD_LOGIC_VECTOR(NB_LANES*3-1 downto 0);
            Xdata: in STD_LOGIC_VECTOR(NB_LANES*XLEN-1 downto 0); --data from scalar register
            Vdata: in STD_LOGIC_VECTOR(2*NB_LANES*64-1 downto 0); --data coming from Register File, 2 since we always have 2 operands
            Idata: in STD_LOGIC_VECTOR(NB_LANES*5-1 downto 0); --data coming from immediate field of size 5 bits
            op1_src: in STD_LOGIC_VECTOR(2*NB_LANES-1 downto 0); -- selects between scalar/vector reg or immediate from operand 2 
                                                -- 00 = vector reg
                                                -- 01 = scalar reg
                                                -- 10 = immediate
                                                -- 11 = RESERVED (unbound)
            funct6: in STD_LOGIC_VECTOR(NB_LANES*6-1 downto 0); --to know which operation
            funct3: in STD_LOGIC_VECTOR (NB_LANES*3-1 downto 0); --to know which operation
            WriteEn_i: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --WriteEn from controller
            WriteEn_o: out STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --WriteEn out to Register File
            WriteEnSel_i: in STD_LOGIC_VECTOR(NB_LANES*8-1 downto 0); --WriteEnSel from OffsetGen
            WriteEnSel_o: out STD_LOGIC_VECTOR(NB_LANES*8-1 downto 0); --WriteEnSel out to Register File
            WriteDest_i : in STD_LOGIC_VECTOR (NB_LANES*(4-(lgNB_LANES-1))-1 downto 0);  
            WriteDest_o : out STD_LOGIC_VECTOR (NB_LANES*(4-(lgNB_LANES-1))-1 downto 0); 
            result: out STD_LOGIC_VECTOR(NB_LANES*64-1 downto 0); --result vector
            w_offset_in : in STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);--write offset coming from offset_generator into EX pipeline reg
            w_offset_out : out STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);--; --write offset coming from WB pipeline reg
            i_done : in STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --coming from offset gen, used to flush control signals of a specific lane
            --done_i: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --done flag coming from offset gen to be rippled through pipeline regs
            o_done: out STD_LOGIC_VECTOR(NB_LANES-1 downto 0) --done flag generated by offset gen coming from WB pipeline reg
            );
end component;

 signal clk:  STD_LOGIC; 
 signal rst:  STD_LOGIC;
 signal mask_reg: STD_LOGIC_VECTOR(VLEN-1 downto 0);
 signal vm:  STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
 signal Xdata:  STD_LOGIC_VECTOR(NB_LANES*XLEN-1 downto 0); --data from scalar register
 signal Vdata:  STD_LOGIC_VECTOR(2*NB_LANES*ELEN-1 downto 0); --data coming from Register File, 2 since we always have 2 operands
 signal Idata:  STD_LOGIC_VECTOR(NB_LANES*5-1 downto 0); --data coming from immediate field of size 5 bits
 signal op1_src:  STD_LOGIC_VECTOR(2*NB_LANES-1 downto 0); -- selects between scalar/vector reg or immediate from operand 2 
 signal funct6:  STD_LOGIC_VECTOR(NB_LANES*6-1 downto 0); --to know which operation
  signal sew:  STD_LOGIC_VECTOR (NB_LANES*3-1 downto 0);
 signal funct3:  STD_LOGIC_VECTOR (NB_LANES*3-1 downto 0); --to know which operation
 signal WriteEn_i:  STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --WriteEn from controller
 signal WriteEn_o:  STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --WriteEn out to Register File
 signal WriteDest_i :  STD_LOGIC_VECTOR (NB_LANES*(4-(lgNB_LANES-1))-1 downto 0);  
 signal WriteDest_o :  STD_LOGIC_VECTOR (NB_LANES*(4-(lgNB_LANES-1))-1 downto 0); 
 signal result:  STD_LOGIC_VECTOR(NB_LANES*ELEN-1 downto 0); --result vector
 signal w_offset_in :  STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);--write offset coming from offset_generator into EX pipeline reg
 signal w_offset_out :  STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);--; --write offset coming from WB pipeline reg
 signal i_done :  STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
 signal  WriteEnSel_i: STD_LOGIC_VECTOR(NB_LANES*8-1 downto 0); --WriteEnSel from OffsetGen
 signal  WriteEnSel_o: STD_LOGIC_VECTOR(NB_LANES*8-1 downto 0); --WriteEnSel to RegFile
begin
    DUT: ALU_with_pipeline --generic map(NB_LANES,VLMAX, ELEN, lgSEW_MAX, XLEN, VLEN)
                           port map(
                         clk          => clk          ,        
                         rst          => rst          ,        
                         mask_reg      => mask_reg    ,    
                         vm           => vm           ,  
                         sew          => sew          ,
                         Xdata        => Xdata        ,      
                         Vdata        => Vdata        ,      
                         Idata        => Idata        ,      
                         op1_src      => op1_src      ,    
                         funct6       => funct6       ,     
                         funct3       => funct3       ,     
                         WriteEn_i    => WriteEn_i    ,
                         WriteEnSel_i => WriteEnSel_i , 
                         WriteEnSel_o => WriteEnSel_o ,
                         WriteEn_o    => WriteEn_o    ,
                         WriteDest_i  => WriteDest_i  , 
                         WriteDest_o  => WriteDest_o  , 
                         result       => result       ,      
                         w_offset_in  => w_offset_in  ,
                         w_offset_out => w_offset_out ,
                         i_done       => i_done     
                           );
                                    
    clk_proc: process begin
        clk<='0';
        wait for 5ns;
        clk<='1'; 
        wait for 5ns;
    end process;
    
    process begin
        rst<='1'; wait for 5ns; rst<= '0'; wait for 5ns;rst<='1';wait for 5ns;
        
        --For testbenching purposes, change ELEN to 32 bits instead of 1024
        
        
        -- Add instruction that adds operands from Vdata since op1_src is 00
        -- Expected result: Lane 0: 5 and Lane 1: 10
        mask_reg<=(others=>'1');
        sew<="000000";
        funct3<= "000000";
        Xdata<= x"0000000600000003";
        Vdata<=x"0202020202020202020202020202020202020202020202020202020202020202";     
        Idata<= "0001100111";
        op1_src<= "0000";
        funct6<="000000000000";
        WriteEn_i<= "11";
        WriteDest_i<="00000000";
        WriteEnSel_i<="0000111100001111";
        vm<="11";
        w_offset_in<="0000000000000001";
        wait for 10ns;
        w_offset_in<="0000000000000000";
        Vdata<=x"0303030303030303030303030320303030303030303030303030303030303030";
        wait for 10ns;
        w_offset_in<="0000000000000001";
        Vdata<=x"0202020202020202020202020202020202020202020202020202020202020202";
        i_done<="11";
       
        wait;
    end process;

end ALU_with_pipeline_tb_arch;
