library IEEE;
library work;
use work.custom_types.all;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity ALU_with_pipeline is
    Port (  clk: in STD_LOGIC; 
            rst: in STD_LOGIC;
            mask_reg: in STD_LOGIC_VECTOR(VLEN-1 downto 0);
            vm: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
            sew: in STD_LOGIC_VECTOR(NB_LANES*3-1 downto 0);
            Xdata: in STD_LOGIC_VECTOR(NB_LANES*XLEN-1 downto 0); --data from scalar register
            Vdata: in STD_LOGIC_VECTOR(2*NB_LANES*64-1 downto 0); --data coming from Register File, 2 since we always have 2 operands
            Idata: in STD_LOGIC_VECTOR(NB_LANES*5-1 downto 0); --data coming from immediate field of size 5 bits
            op1_src: in STD_LOGIC_VECTOR(2*NB_LANES-1 downto 0); -- selects between scalar/vector reg or immediate from operand 2 
                                                -- 00 = vector reg
                                                -- 01 = scalar reg
                                                -- 10 = immediate
                                                -- 11 = RESERVED (unbound)
            funct6: in STD_LOGIC_VECTOR(NB_LANES*6-1 downto 0); --to know which operation
            funct3: in STD_LOGIC_VECTOR (NB_LANES*3-1 downto 0); --to know which operation
            WriteEn_i: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --WriteEn from controller
            WriteEn_o: out STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --WriteEn out to Register File
            WriteEnSel_i: in STD_LOGIC_VECTOR(NB_LANES*8-1 downto 0); --WriteEnSel from OffsetGen
            WriteEnSel_o: out STD_LOGIC_VECTOR(NB_LANES*8-1 downto 0); --WriteEnSel out to Register File
            WriteDest_i : in STD_LOGIC_VECTOR (NB_LANES*(4-(lgNB_LANES-1))-1 downto 0);  
            WriteDest_o : out STD_LOGIC_VECTOR (NB_LANES*(4-(lgNB_LANES-1))-1 downto 0); 
            result: out STD_LOGIC_VECTOR(NB_LANES*64-1 downto 0); --result vector
            w_offset_in : in STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);--write offset coming from offset_generator into EX pipeline reg
            w_offset_out : out STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);--; --write offset coming from WB pipeline reg
            i_done : in STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --coming from offset gen, used to flush control signals of a specific lane
            --done_i: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --done flag coming from offset gen to be rippled through pipeline regs
            o_done: out STD_LOGIC_VECTOR(NB_LANES-1 downto 0) --done flag generated by offset gen coming from WB pipeline reg
            );
end ALU_with_pipeline;

architecture Behavioral of ALU_with_pipeline is
    
component ALU_lane is
    Port (  
            operand1: in STD_LOGIC_VECTOR(63 downto 0);
            operand2: in STD_LOGIC_VECTOR(63 downto 0);
            funct6: in STD_LOGIC_VECTOR (5 downto 0); --to know which operation
            funct3: in STD_LOGIC_VECTOR (2 downto 0); 
            sew: in STD_LOGIC_VECTOR(2 downto 0);
            result: out STD_LOGIC_VECTOR(63 downto 0) 
            );
end component;

component MV_Block is
    Port (  vs1_data: in STD_LOGIC_VECTOR(63 downto 0); -- data from VS1 vector register
            vs2_data: in STD_LOGIC_VECTOR(63 downto 0); -- data from VS2 vector register
            mask_reg: in STD_LOGIC_VECTOR(VLEN-1 downto 0); --mask bit of ith element
            vm: in STD_LOGIC;
            data_out: out STD_LOGIC_VECTOR(ELEN-1 downto 0)
     );
end component;

signal s_operand1: STD_LOGIC_VECTOR(NB_LANES*ELEN-1 downto 0); --Op2 vector (output from mux)

--outputs from pipeline register between RegFile and ALU
signal  s_Xdata:  STD_LOGIC_VECTOR(NB_LANES*XLEN-1 downto 0); --data from scalar register
signal  s_Vdata: STD_LOGIC_VECTOR(2*NB_LANES*64-1 downto 0); --data coming from Register File, 2 since we always have 2 operands
signal  s_Idata:  STD_LOGIC_VECTOR(NB_LANES*5-1 downto 0); --data coming from immediate field of size 5 bits
signal  s_op1_src:  STD_LOGIC_VECTOR(2*NB_LANES-1 downto 0); -- selects between scalar/vector reg or immediate from operand 2                                                                                                                           
signal  s_funct6:  STD_LOGIC_VECTOR(NB_LANES*6-1 downto 0); --to know which operation
signal  s_funct3:  STD_LOGIC_VECTOR (NB_LANES*3-1 downto 0); --to know which operation
signal  s_sew:  STD_LOGIC_VECTOR (NB_LANES*3-1 downto 0);
signal  s_WriteEn_i:  STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --WriteEn from controller
signal  s_WriteDest_i : STD_LOGIC_VECTOR (NB_LANES*(4-(lgNB_LANES-1))-1 downto 0);  
signal  s_vm:  STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
signal  s_w_offset_in :  STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);--offset coming from the pipeline
signal  s_i_done: STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
signal  s_mask_reg: STD_LOGIC_VECTOR(VLEN-1 downto 0);

--signal s_done :  STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --offset going to pipeline
--output from ALU to pipeline register between ALU and WB stage
signal  s_result: STD_LOGIC_VECTOR(NB_LANES*64-1 downto 0); --result vector
signal  s_result_pipeline: STD_LOGIC_VECTOR(NB_LANES*64-1 downto 0); --result vector
signal  a_result: STD_LOGIC_VECTOR(NB_LANES*64-1 downto 0); --result from ALU Lanes
signal  mv_result: STD_LOGIC_VECTOR(NB_LANES*64-1 downto 0); --result from MV Blocks
begin

    pipeline_regs: process(clk, rst,Vdata,Idata,Xdata,op1_src,funct6,funct3,WriteEn_i,WriteEnSel_i,w_offset_in,mask_reg) 
    begin
        if(rst='0') then --reset outputs of pipeline registers
            s_Xdata<=  (others=>'0');
            --s_Vdata<= (others=>'0');
            s_Idata<=  (others=>'0');
            s_op1_src<=(others=>'0');
            s_funct6<= (others=>'0');
            s_funct3<= (others=>'0');    
            result<= (others=>'0');
            s_WriteEn_i<=(others=>'0');
            WriteEn_o<=(others=>'0');
            s_w_offset_in<=(others=>'0');
            --s_done<=(others=>'0');
            w_offset_out<=(others=>'0');
            s_mask_reg<=(others=>'0');
            WriteEnSel_o<=(others=>'0');
            s_WriteDest_i<=(others=>'0');
            
        elsif(rising_edge(clk)) then 
            --s_Vdata<=Vdata;
            s_Xdata<=  Xdata;
            s_Idata<=  Idata; 
            s_mask_reg<=mask_reg;
            s_vm<= vm;
            s_op1_src<=op1_src;
            s_funct6<= funct6;
            s_funct3<= funct3;   
                   
            s_WriteEn_i<=WriteEn_i;
            WriteEn_o<=s_WriteEn_i;
            

            result<=s_result;
            
            
            
            s_WriteDest_i<=WriteDest_i;
            WriteDest_o<=s_WriteDest_i;
            


            --Everything coming from OffsetGen doesn't need another signal
            o_done<=i_done;
            
            w_offset_out<=w_offset_in;
            WriteEnSel_o<=WriteEnSel_i;            
--            s_WriteEnSel_i<=WriteEnSel_i;
--            WriteEnSel_o<=s_WriteEnSel_i;    
--          END_INST: for i in 0 to NB_LANES-1 loop
--            if(i_done(i)='1' and WriteEnSel_i(8*(i+1) downto 8*i)="00000000") then 
--                --busy_lanes(i)<= '0';
--                --vstart(lgVLEN*(i+1)-1 downto lgVLEN*i)<=(others=>'0');                 
--                WriteEn_o(i)<='0';   
--                s_WriteEn_i(i)<='0';
--            end if;
--        end loop;
            
            s_sew<=sew;         
        end if;       
 
    end process;
    
    LANES_GEN:for i in 0 to NB_LANES-1 generate   
    ALU: ALU_lane 
                  port map(
                  operand1=> s_operand1((i+1)*64-1 downto i*64), -- RegFile output is of the form [...Op2,Op1]
                  operand2=>Vdata((2*i+2)*64-1 downto (2*i+1)*64),
                  funct6=> s_funct6((i+1)*6-1 downto i*6),
                  funct3=> s_funct3((i+1)*3-1 downto i*3),
                  sew=> s_sew((i+1)*3-1 downto i*3),
                  result=> a_result((i+1)*64-1 downto i*64)
                    );
    MV: MV_Block  
                  port map(
                  vs1_data=> s_operand1((i+1)*ELEN-1 downto i*ELEN), -- RegFile output is of the form [...Op2,Op1]
                  vs2_data=> Vdata((2*i+2)*ELEN-1 downto (2*i+1)*ELEN),
                  mask_reg=> s_mask_reg,
                  vm=> vm(i),
                  data_out=> mv_result((i+1)*ELEN-1 downto i*ELEN)
                  );

    end generate LANES_GEN;
    
    op2_mux:process(s_op1_src,Vdata,s_Xdata,s_Idata,s_funct6,a_result,mv_result) -- process to select operand2 based on s_op2_src
    begin 
       for i in 0 to NB_LANES-1 loop
            if (s_op1_src(2*i+1 downto 2*i)="00") then
                s_operand1((i+1)*64-1 downto i*64)<=Vdata((2*i+1)*64-1 downto 2*i*64);
            elsif (s_op1_src(2*i+1 downto 2*i)="01") then
                s_operand1((i+1)*64-1 downto i*64)<=std_logic_vector(resize(signed(s_Xdata((i+1)*XLEN-1 downto i*XLEN)),64));--need to sign-extend because XLEN not necessarily = SEW
            elsif (s_op1_src(2*i+1 downto 2*i)="10") then
                s_operand1((i+1)*64-1 downto i*64)<= std_logic_vector(resize(signed(s_Idata((i+1)*5-1 downto i*5)),64));--need to sign-extend because imm is 5 bits
            else 
                s_operand1((i+1)*64-1 downto i*64)<=(others=>'0');
            end if;
            if (s_funct6((i+1)*6-1 downto i*6)="010111") then  
                s_result((i+1)*64-1 downto i*64)<=mv_result((i+1)*64-1 downto i*64);
            else
                s_result((i+1)*64-1 downto i*64)<=a_result((i+1)*64-1 downto i*64);    
            end if;        
        end loop;
   end process;               
end Behavioral;