library IEEE;
library work;
use work.custom_types.all;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity RegFile_ALU is
    Port(   clk: in STD_LOGIC; 
            rst: in STD_LOGIC;
            Xdata: in STD_LOGIC_VECTOR(NB_LANES*XLEN-1 downto 0); --data from scalar register
            Idata: in STD_LOGIC_VECTOR(NB_LANES*5-1 downto 0); --data coming from immediate field of size 5 bits
            op1_src: in STD_LOGIC_VECTOR(2*NB_LANES-1 downto 0); -- selects between scalar/vector reg or immediate from operand 2 
                                                -- 00 = vector reg
                                                -- 01 = scalar reg
                                                -- 10 = immediate
                                                -- 11 = RESERVED (unbound)
            funct6: in STD_LOGIC_VECTOR(NB_LANES*6-1 downto 0); --to know which operation
            funct3: in STD_LOGIC_VECTOR (NB_LANES*3-1 downto 0); --to know which operation
            WriteEn_i: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --WriteEn from controller
            ------Register File            
            sew: in STD_LOGIC_VECTOR (3*NB_LANES-1 downto 0);
            vlmul: in STD_LOGIC_VECTOR(3*NB_LANES-1 downto 0);
            vm: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0);            
            vl: in STD_LOGIC_VECTOR(NB_LANES*XLEN-1 downto 0);
            vstart: in STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);
            newInst: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
            RegSel: in STD_LOGIC_VECTOR((READ_PORTS_PER_LANE*NB_LANES*REGS_PER_BANK)-1 downto 0); 
            WriteDest : in STD_LOGIC_VECTOR (NB_LANES*REGS_PER_BANK-1 downto 0);
            o_done : out STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --going to controller
            reg_out_1: out STD_LOGIC_VECTOR(VLEN-1 downto 0);  --for testing in software 
            reg_out_2: out STD_LOGIC_VECTOR(VLEN-1 downto 0) --for testing in software 
);
end RegFile_ALU;

architecture Structural of RegFile_ALU is

component ALU_with_pipeline is
    Port (  clk: in STD_LOGIC; 
            rst: in STD_LOGIC;
            mask_reg: in STD_LOGIC_VECTOR(VLEN-1 downto 0);
            vm: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
            sew: in STD_LOGIC_VECTOR(NB_LANES*3-1 downto 0);
            Xdata: in STD_LOGIC_VECTOR(NB_LANES*XLEN-1 downto 0); --data from scalar register
            Vdata: in STD_LOGIC_VECTOR(2*NB_LANES*64-1 downto 0); --data coming from Register File, 2 since we always have 2 operands
            Idata: in STD_LOGIC_VECTOR(NB_LANES*5-1 downto 0); --data coming from immediate field of size 5 bits
            op1_src: in STD_LOGIC_VECTOR(2*NB_LANES-1 downto 0); -- selects between scalar/vector reg or immediate from operand 2 
                                                -- 00 = vector reg
                                                -- 01 = scalar reg
                                                -- 10 = immediate
                                                -- 11 = RESERVED (unbound)
            funct6: in STD_LOGIC_VECTOR(NB_LANES*6-1 downto 0); --to know which operation
            funct3: in STD_LOGIC_VECTOR (NB_LANES*3-1 downto 0); --to know which operation
            WriteEn_i: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --WriteEn from controller
            WriteEn_o: out STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --WriteEn out to Register File
            WriteEnSel_i: in STD_LOGIC_VECTOR(NB_LANES*8-1 downto 0); --WriteEnSel from OffsetGen
            WriteEnSel_o: out STD_LOGIC_VECTOR(NB_LANES*8-1 downto 0); --WriteEnSel out to Register File
            WriteDest_i : in STD_LOGIC_VECTOR (NB_LANES*(4-(lgNB_LANES-1))-1 downto 0);  
            WriteDest_o : out STD_LOGIC_VECTOR (NB_LANES*(4-(lgNB_LANES-1))-1 downto 0); 
            result: out STD_LOGIC_VECTOR(NB_LANES*64-1 downto 0); --result vector
            w_offset_in : in STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);--write offset coming from offset_generator into EX pipeline reg
            w_offset_out : out STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);--; --write offset coming from WB pipeline reg
            i_done : in STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --coming from offset gen, used to flush control signals of a specific lane
            --done_i: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --done flag coming from offset gen to be rippled through pipeline regs
            o_done: out STD_LOGIC_VECTOR(NB_LANES-1 downto 0) --done flag generated by offset gen coming from WB pipeline reg
            );
end component;

component RegFile_OffsetGen is
    Port (
            i_clk : in std_logic;
            i_rst: in std_logic;
            newInst: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
            sew: in std_logic_vector (3*NB_LANES-1 downto 0);
            vm: in STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
            vstart: in STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);
            vlmul: in STD_LOGIC_VECTOR(3*NB_LANES-1 downto 0);             
            o_done : out STD_LOGIC_VECTOR(NB_LANES-1 downto 0); 
            mask_bit: out STD_LOGIC;
            OutPort: out STD_LOGIC_VECTOR((READ_PORTS_PER_LANE*NB_LANES*64)-1 downto 0);
            RegSel: in STD_LOGIC_VECTOR((READ_PORTS_PER_LANE*NB_LANES*REGS_PER_BANK)-1 downto 0); 
            WriteEn : in STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
            WriteEnSel_in: in STD_LOGIC_VECTOR(NB_LANES*8-1 downto 0);
            WriteEnSel_out: out STD_LOGIC_VECTOR(NB_LANES*8-1 downto 0);
            WriteData : in STD_LOGIC_VECTOR (NB_LANES*64-1 downto 0);
            WriteDest : in STD_LOGIC_VECTOR (NB_LANES*REGS_PER_BANK-1 downto 0);
            w_offset_in : in STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);--offset coming from the pipeline
            w_offset_out : out STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0); --offset going to pipeline
            vl: in STD_LOGIC_VECTOR(NB_LANES*XLEN-1 downto 0);
            reg_out_1: out STD_LOGIC_VECTOR(VLEN-1 downto 0);  --for testing in software 
            reg_out_2: out STD_LOGIC_VECTOR(VLEN-1 downto 0) --for testing in software   
  );
end component;

signal     s_RegSel: STD_LOGIC_VECTOR((READ_PORTS_PER_LANE*NB_LANES*REGS_PER_BANK)-1 downto 0); 
signal     s_OutPort: STD_LOGIC_VECTOR((READ_PORTS_PER_LANE*NB_LANES*64)-1 downto 0);
signal     s_WriteEn_o: STD_LOGIC_VECTOR(NB_LANES-1 downto 0);
signal     s_result: STD_LOGIC_VECTOR(NB_LANES*ELEN-1 downto 0);
signal     s_mask_bit: STD_LOGIC;
signal     s_mask_reg: STD_LOGIC_VECTOR(VLEN-1 downto 0);
signal     w_offset_in_sig :  STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);--offset coming from the pipeline
signal     w_offset_out_sig :  STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0); --offset going to pipeline
signal     s_done : STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --coming from offset gen
signal     s_o_done : STD_LOGIC_VECTOR(NB_LANES-1 downto 0); --coming from offset gen
signal      s_WriteDest :  STD_LOGIC_VECTOR (NB_LANES*REGS_PER_BANK-1 downto 0);
signal      s_w_offset_in :  STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0);--offset coming from the pipeline
signal      s_w_offset_out :  STD_LOGIC_VECTOR(NB_LANES*lgVLEN-1 downto 0); 


signal s_WriteEnSel_in: STD_LOGIC_VECTOR(NB_LANES*8-1 downto 0);
signal s_WriteEnSel_out: STD_LOGIC_VECTOR(NB_LANES*8-1 downto 0);
begin
-- This process is to pipeline RegSel to allign with its correct offset values
process(clk,RegSel)
begin
    if rising_edge(clk) then
      s_RegSel<=RegSel;  
    end if;
end process;

RF: RegFile_OffsetGen 
           PORT MAP(
           i_clk=>clk,
           i_rst=>rst,
           newInst=>newInst,
           sew=>sew,
           vm=>vm,
           vstart=>vstart,
           vlmul=>vlmul,
           o_done=>s_done,
           mask_bit=>s_mask_bit,
           OutPort=>s_OutPort,
--           RegSel=>RegSel,
           RegSel=>s_RegSel,
           WriteEn=>s_WriteEn_o,
           WriteEnSel_in=> s_WriteEnSel_in,
           WriteEnSel_out=> s_WriteEnSel_out,
           WriteData=>s_result,
           WriteDest=>s_WriteDest,
           w_offset_in=>s_w_offset_in,
           w_offset_out=>s_w_offset_out,
           vl=>vl,
           reg_out_1=>reg_out_1,
           reg_out_2=>reg_out_2
           );
    
ALU: ALU_with_pipeline 
                           port map(
                           clk=>clk,
                           rst=>rst,
                           mask_reg=>s_mask_reg,
                           vm=>vm,
                           sew=>sew,
                           Xdata=>Xdata,
                           Vdata=>s_OutPort,
                           Idata=>Idata, 
                           op1_src=>op1_src,
                           funct6=>funct6,
                           funct3=>funct3,
                           WriteEn_i=>WriteEn_i,
                           WriteEn_o=>s_WriteEn_o,
                           WriteEnSel_i=>s_WriteEnSel_out,
                           WriteEnSel_o=>s_WriteEnSel_in, 
                           WriteDest_i=>WriteDest,
                           WriteDest_o=>s_WriteDest,
                           result=>s_result,
                           w_offset_in=>s_w_offset_out,
                           w_offset_out=>s_w_offset_in,
                           i_done=>s_done,
                           o_done=>s_o_done
                           );

 o_done<=s_o_done;
 
 
end Structural;